-------------------------------------------------------------------------------
--
-- Project					: VGA_ColorBar
-- File name				: VGA_ColorBar.vhd
-- Title					: VGA display test colors
-- Description				:  
--							: 
-- Design library			: N/A
-- Analysis Dependency		: VGA_SYNC.vhd
-- Simulator(s)				: ModelSim-Altera version 6.1g
-- Initialization			: none
-- Notes					: This model is designed for synthesis
--							: Compile with VHDL'93
--
-------------------------------------------------------------------------------
--
-- Revisions
--			Date				Author				Revision		Comments
--		3/11/2008		W.H.Robinson			Rev A			Creation
--		3/13/2012		W.H.Robinson			Rev B			Update for DE2-115 Board
--	  10/31/2014	T. Bruns/M. Beccani		Rev C			Modified to produce rows of colors
--			
-------------------------------------------------------------------------------

-- Always specify the IEEE library in your design
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.all;
USE ieee.std_logic_unsigned.ALL;

-- Entity declaration
ENTITY VGA_ColorBar IS


	PORT
	(
    -- Clocks
    
    CLOCK_50	: IN STD_LOGIC;  -- 50 MHz
 
    -- Buttons 
    
    KEY 		: IN STD_LOGIC_VECTOR (3 downto 0); -- Push buttons

    -- Input switches
    
    SW 			: IN STD_LOGIC_VECTOR (17 downto 0); -- DPDT switches

    -- VGA output
    
    VGA_BLANK_N : out std_logic;            -- BLANK
    VGA_CLK 	 : out std_logic;            -- Clock
    VGA_HS 		 : out std_logic;            -- H_SYNC
    VGA_SYNC_N  : out std_logic;            -- SYNC
    VGA_VS 		 : out std_logic;            -- V_SYNC
    VGA_R 		 : out unsigned(7 downto 0); -- Red[9:0]
    VGA_G 		 : out unsigned(7 downto 0); -- Green[9:0]
    VGA_B 		 : out unsigned(7 downto 0)  -- Blue[9:0]



	);
END VGA_ColorBar;


-- Architecture body 

ARCHITECTURE structural OF VGA_ColorBar IS

COMPONENT VGA_SYNC_module

	PORT(	clock_50Mhz, red, green, blue		: IN	STD_LOGIC;
			red_out, green_out, blue_out, horiz_sync_out, 
			vert_sync_out, video_on, pixel_clock	: OUT	STD_LOGIC;
			pixel_row, pixel_column: OUT STD_LOGIC_VECTOR(9 DOWNTO 0));

END COMPONENT;


SIGNAL red_int				: STD_LOGIC;
SIGNAL green_int	  		: STD_LOGIC;
SIGNAL blue_int     		: STD_LOGIC;
SIGNAL video_on_int		: STD_LOGIC; 
SIGNAL pixel_clock_int	: STD_LOGIC;
SIGNAL pixel_row_int 	: STD_LOGIC_VECTOR(9 DOWNTO 0); 
SIGNAL pixel_column_int : STD_LOGIC_VECTOR(9 DOWNTO 0); 


BEGIN

	VGA_R(6 DOWNTO 0) <= "0000000";
	VGA_G(6 DOWNTO 0) <= "0000000";
	VGA_B(6 DOWNTO 0) <= "0000000";

	U1: VGA_SYNC_module PORT MAP
		(clock_50Mhz		=>	CLOCK_50,
		 red					=>	pixel_row_int(7),
		 green				=>	pixel_row_int(6),	
		 blue					=>	pixel_row_int(5),
		 red_out				=>	VGA_R(7),
		 green_out			=>	VGA_G(7),
		 blue_out			=>	VGA_B(7),
		 horiz_sync_out	=>	VGA_HS,
		 vert_sync_out		=>	VGA_VS,
		 video_on			=>	VGA_BLANK_N,
		 pixel_clock		=>	VGA_CLK,
		 pixel_row			=>	pixel_row_int,
		 pixel_column		=>	pixel_column_int
		);

END structural;

