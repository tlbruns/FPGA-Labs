
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity top_level is
    Port ( CLOCK_50          : in  STD_LOGIC;
           
			  GPIO : inout std_logic_vector(35 downto 0);
           config_finished : out STD_LOGIC;
         --  vga_r     : out  STD_LOGIC_vector(2 downto 0);
         --  vga_g     : out  STD_LOGIC_vector(2 downto 0);
          -- vga_b     : out  STD_LOGIC_vector(2 downto 1);
           

		
--		OV7670_SIOC  : out   STD_LOGIC;
--		OV7670_SIOD  : inout STD_LOGIC;
--		OV7670_RESET : out   STD_LOGIC;
--		OV7670_PWDN  : out   STD_LOGIC;
--		OV7670_VSYNC : in    STD_LOGIC;
--		OV7670_HREF  : in    STD_LOGIC;
--		OV7670_PCLK  : in    STD_LOGIC;
--		OV7670_XCLK  : out   STD_LOGIC;
--		OV7670_D     : in    STD_LOGIC_VECTOR(7 downto 0);

	--	LEDG         : out    STD_LOGIC_VECTOR(7 downto 0);
		
		VGA_HS  		 : out  STD_LOGIC;  -- H_SYNC
		VGA_VS 		 : out  STD_LOGIC;  -- V_SYNC
		VGA_BLANK_N  : out std_logic;   -- BLANK
		VGA_CLK 	 	 : out std_logic;   -- Clock
		VGA_SYNC_N   : out std_logic;   -- SYNC

		VGA_R     	 : out   STD_LOGIC_VECTOR(7 downto 0);
		VGA_G    	 : out   STD_LOGIC_VECTOR(7 downto 0);
		VGA_B        : out   STD_LOGIC_VECTOR(7 downto 0);
		
		KEY 		    : in    STD_LOGIC_VECTOR(3 downto 0)
			  		  
           );
end top_level;

architecture Behavioral of top_level is

	COMPONENT VGA
	PORT(
		CLK25 : IN std_logic;    
		Hsync : OUT std_logic;
		Vsync : OUT std_logic;
		Nblank : OUT std_logic;      
		clkout : OUT std_logic;
		activeArea : OUT std_logic;
		Nsync : OUT std_logic
		);
	END COMPONENT;

	COMPONENT ov7670_controller
	PORT(
		clk : IN std_logic;
		resend : IN std_logic;    
		siod : INOUT std_logic;      
		config_finished : OUT std_logic;
		sioc : OUT std_logic;
		reset : OUT std_logic;
		pwdn : OUT std_logic;
		xclk : OUT std_logic
		);
	END COMPONENT;

	COMPONENT debounce
	PORT(
		clk : IN std_logic;
		i : IN std_logic;          
		o : OUT std_logic
		);
	END COMPONENT;

	COMPONENT frame_buffer
	PORT(
		data : IN std_logic_vector(11 downto 0);
		rdaddress : IN std_logic_vector(16 downto 0);
		rdclock : IN std_logic;
		wraddress : IN std_logic_vector(16 downto 0);
		wrclock : IN std_logic;
		wren : IN std_logic;          
		q : OUT std_logic_vector(11 downto 0)
		);
	END COMPONENT;
	

	COMPONENT ov7670_capture
	PORT(
		pclk : IN std_logic;
		vsync : IN std_logic;
		href : IN std_logic;
		d : IN std_logic_vector(7 downto 0);          
		addr : OUT std_logic_vector(18 downto 0);
		dout : OUT std_logic_vector(11 downto 0);
		we : OUT std_logic
		);
	END COMPONENT;

	COMPONENT RGB
	PORT(
		Din : IN std_logic_vector(11 downto 0);
		Nblank : IN std_logic;          
		R : OUT std_logic_vector(7 downto 0);
		G : OUT std_logic_vector(7 downto 0);
		B : OUT std_logic_vector(7 downto 0)
		);
	END COMPONENT;

	COMPONENT vga_pll
	PORT(
		inclk0 : IN std_logic;          
		c0 : OUT std_logic;
		c1 : OUT std_logic
		);
	END COMPONENT;


	COMPONENT Adress_Generator
	PORT(
		CLK25 : IN std_logic;
		enable : IN std_logic;       
      vsync  : in  	STD_LOGIC;
		adress : INOUT std_logic_vector(16 downto 0)
		);
	END COMPONENT;



   signal clk_camera : std_logic;
   signal clk_vga    : std_logic;
   signal wren       : std_logic;
   signal resend     : std_logic;
   signal nBlank     : std_logic;
   signal vsync      : std_logic;
   signal nSync      : std_logic;
   
   signal wraddress  : std_logic_vector(18 downto 0);
   signal wrdata     : std_logic_vector(11 downto 0);
   signal rdaddress  : std_logic_vector(16 downto 0);
   signal rddata     : std_logic_vector(11 downto 0);
   signal red,green,blue : std_logic_vector(7 downto 0);
   signal activeArea : std_logic;
	
	
begin
   vga_r <= red(7 downto 0);
   vga_g <= green(7 downto 0);
   vga_b <= blue(7 downto 0);
   
	Inst_vga_pll: vga_pll PORT MAP(
		inclk0 => CLOCK_50,
		c0 => clk_camera,
		c1 => clk_vga
	);

   VGA_VS <= vsync;
   
	Inst_VGA: VGA PORT MAP(
		CLK25      => clk_vga,
		clkout     => VGA_CLK,
		Hsync      => VGA_HS,
		Vsync      => vsync,
		Nblank     => VGA_BLANK_N,
		Nsync      => VGA_SYNC_N,
      activeArea => activeArea
	);

	Inst_debounce: debounce PORT MAP(
		clk => CLOCK_50,
		i   => KEY(0),
		o   => resend
	);

	Inst_ov7670_controller: ov7670_controller PORT MAP(
		clk             => clk_camera,
		resend          => resend,
		config_finished => config_finished,
		sioc            => GPIO(24),--ov7670_sioc,
		siod            => GPIO(25),--ov7670_siod,
		reset           => GPIO(10),--ov7670_reset,
		pwdn            => GPIO(11),--ov7670_pwdn,
		xclk            => GPIO(21)--ov7670_xclk
	);

	Inst_frame_buffer: frame_buffer PORT MAP(
		rdaddress => rdaddress,
		rdclock   => clk_vga,
		q         => rddata,
      
		wrclock   => GPIO(20),--ov7670_pclk,
		wraddress => wraddress(16 downto 0),
		data      => wrdata,
		wren      => wren
	);
   
	Inst_ov7670_capture: ov7670_capture PORT MAP(
		pclk  => GPIO(20),--ov7670_pclk,
		vsync => GPIO(22),--ov7670_vsync,
		href  => GPIO(23),--ov7670_href,
		d     => GPIO(19 downto 12),--ov7670_data,
		addr  => wraddress,
		dout  => wrdata,
		we    => wren
	);

	Inst_RGB: RGB PORT MAP(
		Din => rddata,
		Nblank => activeArea,
		R => red,
		G => green,
		B => blue
	);

	Inst_Adress_Generator: Adress_Generator PORT MAP(
		CLK25 => clk_vga,
		enable => activeArea,
      vsync  => vsync,
		adress => rdaddress
	);

end Behavioral;

