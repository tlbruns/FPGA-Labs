library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity icon_takephoto is
	port( index	:	in	integer range 1 to 2500;
			pixel	:	out std_logic_vector(11 downto 0)
			);
end icon_takephoto;

architecture structural of icon_takephoto is

	type icon_t is array(1 to 2500) of std_logic_vector(11 downto 0);
	constant icon_photo : icon_t := ("000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001000100010",
				"011001100110",
				"100110011001",
				"101110111011",
				"110111011101",
				"111011101110",
				"111111111111",
				"111111111111",
				"111011101110",
				"110111011101",
				"101110111011",
				"100110011001",
				"011001100110",
				"001000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001000100010",
				"100010001000",
				"110011001100",
				"111111111111",
				"110111011101",
				"101110111011",
				"100010001000",
				"011001100110",
				"010101010101",
				"010001000100",
				"010001000100",
				"010101010101",
				"011001100110",
				"100010001000",
				"101110111011",
				"110111011101",
				"111111111111",
				"110011001100",
				"100010001000",
				"001000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001100110011",
				"101010101010",
				"111111111111",
				"110111011101",
				"100010001000",
				"001100110011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001100110011",
				"100010001000",
				"110111011101",
				"111111111111",
				"101010101010",
				"001100110011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"101010101010",
				"111111111111",
				"110011001100",
				"010001000100",
				"000000000000",
				"000000000000",
				"000000000000",
				"010001000100",
				"100010001000",
				"101110111011",
				"110011001100",
				"110111011101",
				"111011101110",
				"111011101110",
				"110111011101",
				"110011001100",
				"101110111011",
				"100010001000",
				"010001000100",
				"000000000000",
				"000000000000",
				"000000000000",
				"010001000100",
				"110011001100",
				"111111111111",
				"101010101010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"010101010101",
				"111011101110",
				"110111011101",
				"010001000100",
				"000000000000",
				"000000000000",
				"010001000100",
				"101010101010",
				"111011101110",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101110",
				"101010101010",
				"010001000100",
				"000000000000",
				"000000000000",
				"010101010101",
				"110111011101",
				"111011101110",
				"010101010101",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"100010001001",
				"111111111111",
				"100010001000",
				"000000000000",
				"000000000000",
				"010101010101",
				"110011001100",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111111111111",
				"111111111111",
				"111111111111",
				"110011001100",
				"010101010101",
				"000000000000",
				"000000000000",
				"100010001000",
				"111111111111",
				"100010001001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"101110111011",
				"111111111111",
				"010001000100",
				"000000000000",
				"000100010001",
				"101110111011",
				"111111111111",
				"111111111111",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111111111111",
				"111111111111",
				"101110111011",
				"000100010001",
				"000000000000",
				"010001000100",
				"111111111111",
				"101110111011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"110011001100",
				"111011101110",
				"001000100010",
				"000000000000",
				"010101010101",
				"111111111111",
				"111111111111",
				"111011101110",
				"111011011110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111111111111",
				"111111111111",
				"010101010101",
				"000000000000",
				"001000100010",
				"111011101110",
				"110011001100",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"101110111011",
				"111011101110",
				"000100010001",
				"000000000000",
				"100010001000",
				"111111111111",
				"111111111111",
				"110111011101",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"110111011101",
				"111111111111",
				"111111111111",
				"100010001000",
				"000000000000",
				"000100010001",
				"111011101110",
				"101110111011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"100110011001",
				"111111111111",
				"001000100010",
				"000000000000",
				"100010001000",
				"111111111111",
				"111011101110",
				"110111011101",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"111011101110",
				"111111111111",
				"100010001000",
				"000000000000",
				"001000100010",
				"111111111111",
				"100110011001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"010001000100",
				"111111111111",
				"010001000100",
				"000000000000",
				"011101110111",
				"111111111111",
				"111011101110",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"111011101110",
				"111111111111",
				"011101110111",
				"000000000000",
				"010001000100",
				"111111111111",
				"010001000100",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"111111111111",
				"011101111000",
				"000000000000",
				"010001000100",
				"111111111111",
				"111011101110",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"111011101110",
				"111111111111",
				"010001000100",
				"000000000000",
				"011101110111",
				"111111111111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"100110011001",
				"110111011101",
				"000000000000",
				"000100010001",
				"111011101110",
				"111011101111",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"111011101111",
				"111011101110",
				"000100010001",
				"000000000000",
				"110111011101",
				"100110011001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001000100010",
				"111111111111",
				"001100110011",
				"000000000000",
				"101010101010",
				"111111111111",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"111111111111",
				"101010101010",
				"000000000000",
				"001100110011",
				"111111111111",
				"001000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"101010101010",
				"101110111011",
				"000000000000",
				"001100110011",
				"111111111111",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"111111111111",
				"001100110011",
				"000000000000",
				"101110111011",
				"101010101010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"111111111111",
				"001100110011",
				"000000000000",
				"101110111011",
				"111111111111",
				"110011001101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110011011101",
				"110111011101",
				"110111011110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"110111011110",
				"110111011101",
				"110011011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110011011101",
				"110011001101",
				"111111111111",
				"101110111011",
				"000000000000",
				"001100110011",
				"111111111111",
				"000100010001",
				"000000000000",
				"000000000000",
				"011101110111",
				"110011001100",
				"000000000000",
				"001000100010",
				"111011101111",
				"110111011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110111011101",
				"111011101110",
				"110011001100",
				"101010101010",
				"101010101010",
				"101010101011",
				"101010101010",
				"101010101010",
				"101010101010",
				"110011001100",
				"111011101110",
				"110111011101",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011001101",
				"110111011101",
				"111011101111",
				"001000100010",
				"000000000000",
				"110011001100",
				"011101110111",
				"000000000000",
				"000000000000",
				"110011001100",
				"011101110111",
				"000000000000",
				"100010001001",
				"111111111111",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001100",
				"110111011110",
				"111011101110",
				"111111111111",
				"111011101110",
				"011101110111",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"011101110111",
				"111011101110",
				"111111111111",
				"111011101110",
				"110111011101",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001101",
				"110011001100",
				"111111111111",
				"100010001001",
				"000000000000",
				"011101110111",
				"110011001100",
				"000000000000",
				"000100010001",
				"111011101110",
				"001000100010",
				"000000000000",
				"110011001100",
				"110111011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111011110",
				"101010111011",
				"011101110111",
				"100010001000",
				"011001100110",
				"000100010001",
				"001000100010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"000100010001",
				"011001100110",
				"100010001000",
				"011101110111",
				"101010111011",
				"110111011110",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111011101",
				"110011001100",
				"000000000000",
				"001000100010",
				"111011101110",
				"000100010001",
				"010101010101",
				"110011001100",
				"000000000000",
				"001000100010",
				"111011101110",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111011101",
				"100110011010",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"001100110011",
				"001100110011",
				"001000100010",
				"001000100010",
				"001100110011",
				"001100110011",
				"001000100010",
				"001000100010",
				"010000110100",
				"001100110100",
				"000100010010",
				"000100010001",
				"000100010001",
				"000100010010",
				"100110011010",
				"110111011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"111011101110",
				"001000100010",
				"000000000000",
				"110011001100",
				"010101010101",
				"100010001000",
				"100110011001",
				"000000000000",
				"011001100110",
				"111011101110",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111011101",
				"010001000100",
				"000100010001",
				"010001000100",
				"001100110100",
				"001100110011",
				"001100110011",
				"001000100010",
				"010101010101",
				"100110011001",
				"101110111011",
				"101110111011",
				"100110011001",
				"010101010101",
				"001000100010",
				"001100110011",
				"001100110011",
				"001100110011",
				"010001000100",
				"000100010001",
				"010001000101",
				"110111011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"111011101110",
				"011001100110",
				"000000000000",
				"100110011001",
				"100010001000",
				"101010101010",
				"011101110111",
				"000000000000",
				"100010001000",
				"111011101110",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"010101010101",
				"001000100010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"011001100110",
				"110111011101",
				"111111111111",
				"111011101110",
				"111011101110",
				"111111111111",
				"110111011101",
				"011001100110",
				"001000100010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"010101010101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"111011101110",
				"100010001000",
				"000000000000",
				"011101110111",
				"101010101010",
				"101110111011",
				"010101010101",
				"000000000000",
				"100110011010",
				"110111011101",
				"101111001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"010101010101",
				"001000100010",
				"001100110011",
				"001100110011",
				"001000100010",
				"010001000101",
				"110111011101",
				"111011011110",
				"100010001000",
				"010001000100",
				"010001000100",
				"100010001000",
				"111011101110",
				"110111011101",
				"010001000101",
				"001000100010",
				"001100110011",
				"001100110011",
				"001000100010",
				"010101010101",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110111011101",
				"100110101010",
				"000000000000",
				"010101010101",
				"101110111011",
				"110011001100",
				"010001000100",
				"000000000000",
				"101010101010",
				"110011001101",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"110011001100",
				"110011001100",
				"010101010101",
				"001000100010",
				"001100110011",
				"001100110011",
				"001000100010",
				"100110011001",
				"111011111111",
				"100010001000",
				"000000000001",
				"000100010001",
				"000100010001",
				"000000000001",
				"100010001000",
				"111111111111",
				"100110011001",
				"001000100010",
				"001100110011",
				"001100110011",
				"001000100010",
				"010101010101",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"110011001101",
				"101010101010",
				"000000000000",
				"010001000100",
				"110011001100",
				"110011001101",
				"001100110011",
				"000000000000",
				"101110111011",
				"110011001100",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"110011001100",
				"010101010101",
				"001000100010",
				"001100110011",
				"001100110011",
				"001100110011",
				"101010111011",
				"110111011101",
				"010001000100",
				"001000100010",
				"001100110011",
				"001100110011",
				"001000100010",
				"010001000100",
				"110111011101",
				"101110111011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"010101010101",
				"110011001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"110011001100",
				"101110111011",
				"000000000000",
				"001100110011",
				"110011001101",
				"110011001100",
				"001100110011",
				"000000000000",
				"101010101011",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"110011001100",
				"010101010101",
				"001000100010",
				"001100110011",
				"001100110011",
				"001100110011",
				"101010101010",
				"110011011101",
				"010001000100",
				"001000100010",
				"001100110011",
				"001100110011",
				"001000100010",
				"010001000100",
				"110111001101",
				"101010101010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"010101010101",
				"110011001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"101010101011",
				"000000000000",
				"001100110011",
				"110011001101",
				"101111001100",
				"010001000100",
				"000000000000",
				"101010101010",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"010101010101",
				"001000100010",
				"001100110011",
				"001100110011",
				"001000100010",
				"100010001000",
				"111011101110",
				"100010001000",
				"000100010001",
				"001000100010",
				"001000100010",
				"000100010001",
				"100010001000",
				"111011101110",
				"100010001000",
				"001000100010",
				"001100110011",
				"001100110011",
				"001000100010",
				"010101010101",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"101010101010",
				"000000000000",
				"010001000100",
				"110010111100",
				"101110111011",
				"010101010101",
				"000000000000",
				"100110011001",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"010001010101",
				"001000100010",
				"001100110011",
				"001100110011",
				"001000100010",
				"010001000100",
				"110011001100",
				"110111011101",
				"100010001000",
				"010001000100",
				"010001000100",
				"100010001000",
				"110111011101",
				"110011001100",
				"010001000100",
				"001000100010",
				"001100110011",
				"001100110011",
				"001000100010",
				"010001010101",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"100110011001",
				"000000000000",
				"010101010101",
				"101110111011",
				"100110011001",
				"011101110111",
				"000000000000",
				"011101111000",
				"110011011101",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"010001000101",
				"001000100010",
				"001100110011",
				"001100110011",
				"001100110011",
				"000100010001",
				"010101010101",
				"110011001100",
				"111011101110",
				"110011001101",
				"110011001101",
				"111011101110",
				"110011001100",
				"010101010101",
				"000100010001",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"010001000101",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001101",
				"011101111000",
				"000000000000",
				"011101110111",
				"100110011001",
				"011101110111",
				"100110011001",
				"000000000000",
				"010101010101",
				"110011011101",
				"101010101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"010001000100",
				"001000100010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"000100010001",
				"010001000100",
				"100010001000",
				"101010101010",
				"101010101010",
				"100010001000",
				"010001000100",
				"000100010001",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"010001000100",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"110011011101",
				"010101010101",
				"000000000000",
				"100110011001",
				"011101110111",
				"010001000100",
				"101010101011",
				"000000000000",
				"001000100010",
				"110011001100",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101110111100",
				"010001000101",
				"000100010001",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"000100010001",
				"001000100010",
				"001000100010",
				"000100010001",
				"001000100010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"000100010001",
				"010001000101",
				"110010111100",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"110011001100",
				"001000100010",
				"000000000000",
				"101010101011",
				"010001000100",
				"000100010001",
				"110011001100",
				"001000100010",
				"000000000000",
				"101010101010",
				"101110111011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101010",
				"101010101011",
				"101010101011",
				"101110111011",
				"100110011001",
				"001100110011",
				"000100010001",
				"000100010001",
				"000100010010",
				"000100010001",
				"000100010001",
				"000100010010",
				"000100010010",
				"000100010001",
				"000100010001",
				"000100010010",
				"000100010010",
				"000100010001",
				"000100010001",
				"000100010010",
				"000100010001",
				"000100010001",
				"001100110011",
				"100110011001",
				"101110111011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101010",
				"101010101010",
				"101010101011",
				"101110111011",
				"101010101010",
				"000000000000",
				"001000100010",
				"110011001100",
				"000100010001",
				"000000000000",
				"101010101010",
				"011001100110",
				"000000000000",
				"011101110111",
				"110011001100",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111100",
				"101010101010",
				"011101111000",
				"100001111000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011101111000",
				"101010101010",
				"101110111100",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"110011001100",
				"011101110111",
				"000000000000",
				"011001100111",
				"101010101010",
				"000000000000",
				"000000000000",
				"010101010101",
				"101010101010",
				"000000000000",
				"001000010001",
				"101111001100",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101111001100",
				"001000100010",
				"000000000000",
				"101010101010",
				"010101010101",
				"000000000000",
				"000000000000",
				"000100010001",
				"110011001100",
				"010000110100",
				"000000000000",
				"100010001000",
				"101110111100",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111100",
				"100010001000",
				"000000000000",
				"001100110100",
				"110011001100",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"011101111000",
				"100110011001",
				"000000000000",
				"001000100010",
				"101111001100",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101111001100",
				"001000100010",
				"000000000000",
				"100110011001",
				"011101111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"110011001100",
				"010001000100",
				"000000000000",
				"011101110111",
				"101110111100",
				"100110011010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110011010",
				"101110111100",
				"011101110111",
				"000000000000",
				"010001000100",
				"110011001100",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"011001100111",
				"101110111011",
				"000000000000",
				"000000000000",
				"101010101010",
				"101010101011",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"101010101011",
				"101010101010",
				"000000000000",
				"000000000000",
				"101010101011",
				"011001100111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"101111001100",
				"011101110111",
				"000000000000",
				"001000100010",
				"101110111011",
				"101010101010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011001",
				"101010101010",
				"101110111011",
				"001000100010",
				"000000000000",
				"011101110111",
				"101110111100",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001100110011",
				"110011001100",
				"010001000100",
				"000000000000",
				"010001000100",
				"101110111100",
				"100110011010",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011010",
				"101110111100",
				"010001000100",
				"000000000000",
				"010001000100",
				"110011001100",
				"001100110011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"011001100110",
				"101110111100",
				"001100110011",
				"000000000000",
				"010101010101",
				"101110111011",
				"100110101010",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110101010",
				"101110111011",
				"010101010101",
				"000000000000",
				"001100110011",
				"101110111100",
				"011001100110",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"011101110111",
				"101110111011",
				"001000100010",
				"000000000000",
				"010001000100",
				"101110111011",
				"101010101010",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101110111011",
				"010001000100",
				"000000000000",
				"001000100010",
				"101110111011",
				"011101111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"100010001000",
				"101110111011",
				"001100110011",
				"000000000000",
				"001000100010",
				"100110011001",
				"101010111011",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101110111011",
				"100110011010",
				"001000100010",
				"000000000000",
				"001100110011",
				"101110111011",
				"100010001000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"011101110111",
				"101110111011",
				"010101010101",
				"000000000000",
				"000000000000",
				"011001100110",
				"101010101010",
				"101010101010",
				"100110011001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"011001100110",
				"000000000000",
				"000000000000",
				"010101010101",
				"101110111011",
				"011101110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"010101010101",
				"101110111100",
				"100010001000",
				"000000000000",
				"000000000000",
				"001000100010",
				"011101110111",
				"101010101010",
				"101010101010",
				"100110011010",
				"100110011001",
				"100010001001",
				"100010001001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010001001",
				"100010001001",
				"100010001001",
				"100010001001",
				"100010001001",
				"100010011001",
				"100110011010",
				"101010101010",
				"101010101010",
				"011101110111",
				"001000100010",
				"000000000000",
				"000000000000",
				"011110001000",
				"101110111100",
				"010101010101",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001100110011",
				"101010101010",
				"101010101010",
				"010101010101",
				"000000000000",
				"000000000000",
				"000100010001",
				"010101010110",
				"100010001000",
				"100110011010",
				"101010101010",
				"101010101010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011001",
				"100110011010",
				"100110011010",
				"101010101010",
				"101010101010",
				"100110011010",
				"100010001000",
				"010101010110",
				"001000100010",
				"000000000000",
				"000000000000",
				"010101010101",
				"101010101010",
				"101010101010",
				"001100110011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"010101010110",
				"101110111011",
				"100110011001",
				"010101010101",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"010001000100",
				"010101010101",
				"011001100111",
				"011101110111",
				"011101111000",
				"011110001000",
				"011101110111",
				"011001100111",
				"010101010101",
				"010001000100",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"010101010101",
				"100110011001",
				"101110111011",
				"010101010110",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"011001100110",
				"101010101011",
				"101010101010",
				"011101110111",
				"010001000100",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"010001000100",
				"011101110111",
				"100110011010",
				"101010101011",
				"011001100110",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"010001000100",
				"100010001000",
				"101010101011",
				"101010101010",
				"100010001001",
				"011101110111",
				"011001100110",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100110",
				"011101110111",
				"100010001001",
				"101010101010",
				"101010101011",
				"100010001000",
				"010001000100",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001100110011",
				"010101010101",
				"011101110111",
				"100010001000",
				"100110011001",
				"101010101010",
				"101010101010",
				"100110011001",
				"100010001000",
				"011101110111",
				"010101010101",
				"001100110011",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000"
				);
				
begin
	pixel <= icon_photo(index);

end structural; 
	
			